LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY cnt4 IS
	PORT(CLK:IN STD_LOGIC;
	 CQ:OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END cnt4;
ARCHITECTURE behav OF cnt4 IS
BEGIN
	PROCESS(CLK)
	 VARIABLE CQI:STD_LOGIC_VECTOR(3 DOWNTO 0);
	BEGIN
	  IF CLK'EVENT AND CLK='1' THEN
		CQI:=CQI+1;
	  END IF;
	CQ<=CQI;
   END PROCESS;
  END behav;
	